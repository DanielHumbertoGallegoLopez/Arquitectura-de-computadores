--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   17:02:03 04/17/2017
-- Design Name:   
-- Module Name:   C:/Users/utp.CRIE/Desktop/Procesador_2_PruebasModulos/Procesador_2/Prueba_sEU.vhd
-- Project Name:  Procesador_2
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: sEU
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY Prueba_sEU IS
END Prueba_sEU;
 
ARCHITECTURE behavior OF Prueba_sEU IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT sEU
    PORT(
         imm13 : IN  std_logic_vector(12 downto 0);
         SalidaSEU : OUT  std_logic_vector(31 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal imm13 : std_logic_vector(12 downto 0) := (others => '0');

 	--Outputs
   signal SalidaSEU : std_logic_vector(31 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: sEU PORT MAP (
          imm13 => imm13,
          SalidaSEU => SalidaSEU
        );
 

   -- Stimulus process
   stim_proc: process
   begin		
      
		imm13 <= "0100111001010";

      wait;
   end process;

END;
